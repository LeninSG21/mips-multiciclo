module data_reg (
        
    );
    

endmodule