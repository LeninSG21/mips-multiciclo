module rf(
  //We are asuming always enabled RAM
  input clk, we, rst,
  input [4:0] rs_add,
  input [4:0] rt_add,
  input [4:0] rd_add,
  input [31:0] rd_data,
  output reg [31:0] rs_data,
  output reg [31:0] rt_data
  );
  
  reg [31:0] mem[31:0];
  int i;
  
  initial
  begin
  	$readmemh("memfile.dat", mem);
  end
  
  always @ (posedge clk or rst)
  begin

      if(rst)
        for(i = 0; i <= 31; i = i+1)
          mem[i] <= 0;
      else if(we)
        begin
          if(rd_add != 0)
            begin
            mem[rd_add] <= rd_data;
            $writememh("memfile2.dat", mem);
            end
        end
  end
 
  assign rs_data = mem[rs_add];
  assign rt_data = mem[rt_add];
  
endmodule
